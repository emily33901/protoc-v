module compiler

// TODO this file needs a massive refactor and clean
// So much code just everywhere with functions that dont
// make any sense
// Please just fix it before its too late...

// Other things that would be nice

// Functions for getting names / types consistently
// instead of manually creating m_name and m_full_name
// in each of the places that they are used!

struct Gen {
	type_table &TypeTable
	w Writer

mut: 
	// Maps proto packages to v packages
	package_lookup map[string]string

	current_package string
}

fn (mut g Gen) gen_file_header(f &File) {
	// TODO figure out an appropriate module
	// if the file doesnt have an explicit package set

	mut mod := ''
	for _, o in f.options {
		if o.ident == 'v_package' {
			mod = o.value.value
		}
	}

	if mod == '' {
		mod = f.package.all_after_last('.')
	}

	g.w.l('
// Generated by vproto - Do not modify
module ${mod}

import emily33901.vproto

')

	for _, i in f.imports {
		x := i.package
		g.w.l('import ${g.package_lookup[x]}')
	}

// g.w.l('
// pub const (
// 	v_package = \'$g.current_package\'
// )')

}

fn (mut g Gen) gen_enum_definition(type_context []string, e &Enum) {
	names := g.message_names(type_context, e.name)
	
	e_name := names.struct_name
	e_full_name := names.lowercase_name

	g.w.l('enum ${e_name} {')

	for _, field in e.fields {
		g.w.l('${to_v_field_name(field.name)} = $field.value.value')
	}

	g.w.l('}')

	// generate packing and unpacking functions

	g.w.l('fn pack_${e_full_name}(e $e_name, num u32) []byte {')
	g.w.l('return vproto.pack_int32_field(int(e), num)')
	g.w.l('}')

	g.w.l('fn unpack_${e_full_name}(buf []byte, tag_wiretype vproto.WireType) (int, $e_name) {')
	g.w.l('i, v := vproto.unpack_int32_field(buf, tag_wiretype)')
	g.w.l('return i, ${e_name}(v)')
	g.w.l('}')

	// TODO helper functions here 
	// https://developers.google.com/protocol-buffers/docs/reference/cpp-generated#enum
}

// TODO When type_to_type changes name change this name too ! 
fn (mut g Gen) type_to_typename(context []string, t string) (string, TypeType) {

	// mut full_context := []string{}
	// full_context << g.current_package.split('.')
	// full_context << context

	return type_to_typename(g.current_package, g.type_table, context, t)
}

fn (g Gen) message_names(context []string, t string) MessageNames {
	return message_names(g.current_package, g.type_table, context, t)
}

fn (g &Gen) type_pack_name(pack_or_unpack string, field_proto_type string, field_v_type string, field_type_type TypeType) string {
	// TODO clean up this whackness :(
	match field_type_type {
		.other {
			match field_proto_type {
				'fixed32' {
					return 'vproto.${pack_or_unpack}_32bit_field'
				}

				'sfixed32' {
					return 'vproto.${pack_or_unpack}_s32bit_field'
				}

				'float' {
					return 'vproto.${pack_or_unpack}_float_field'
				}

				'fixed64' {
					return 'vproto.${pack_or_unpack}_64bit_field'
				}

				'sfixed64' {
					return 'vproto.${pack_or_unpack}_s64bit_field'
				}

				'double' {
					return 'vproto.${pack_or_unpack}_double_field'
				}

				'int32' {
					return 'vproto.${pack_or_unpack}_int32_field'
				}

				'sint32' {
					return 'vproto.${pack_or_unpack}_sint32_field'
				}

				'sint64' {
					return 'vproto.${pack_or_unpack}_sint64_field'
				}

				'uint32' {
					return 'vproto.${pack_or_unpack}_uint32_field'
				}

				'int64' {
					return 'vproto.${pack_or_unpack}_int64_field'
				}

				'uint64' {
					return 'vproto.${pack_or_unpack}_uint64_field'
				}

				'bool' {
					return 'vproto.${pack_or_unpack}_bool_field'
				}

				'string' {
					return 'vproto.${pack_or_unpack}_string_field'
				}

				'bytes' {
					return 'vproto.${pack_or_unpack}_bytes_field'
				}

				else {
					panic('unknown type `$field_proto_type`')
				}
			}
		}

		.enum_, .message {
			return '${pack_or_unpack}_$field_v_type'
		}
	}
}

fn (g &Gen) gen_field_pack_text(
	label, field_proto_type, field_v_type string, 
	field_TypeType TypeType, 
	name, number string, 
	is_packed bool
) (string, string) {
	mut pack_text := ''
	mut unpack_text := ''

	// TODO this isnt ideal

	field_v_type_no_mod := field_v_type.all_after_last('.')
	field_v_type_mod := if field_v_type.contains('.') { field_v_type.all_before_last('.') + '.' } else { '' }

	pack_inside := g.type_pack_name('${field_v_type_mod}pack', field_proto_type, field_v_type_no_mod, field_TypeType)
	unpack_inside := g.type_pack_name('${field_v_type_mod}unpack', field_proto_type, field_v_type_no_mod, field_TypeType)

	match label {
		'optional', 'required' {
			unpack_text += '$number {\n'

			if label == 'optional' {
				pack_text += 'if o.has_$name {\n'

				unpack_text += 'res.has_$name = true\n'
			}

			pack_text += 'res << ${pack_inside}(o.$name, $number)\n'

			if label == 'optional' {
				pack_text += '}\n'
			}

			// unpack text at this point is inside of a match statement checking tag numbers

			// TODO make this into a oneliner again once match bug is fixed

			unpack_text += 'ii, v := ${unpack_inside}(cur_buf, tag_wiretype.wire_type)\n'
			unpack_text += 'res.$name = v\n'
			unpack_text += 'i = ii\n'
			unpack_text += '}\n'
		}
 
		'repeated' {
			if !is_packed {
				pack_text += '// [packed=false]\n'
				pack_text += 'for _, x in o.$name {\n'
				pack_text += 'res << ${pack_inside}(x, $number)\n'
				pack_text += '}\n'

				unpack_text += '$number {\n'
				unpack_text += '// [packed=false]\n'
				unpack_text += 'ii, v := ${unpack_inside}(cur_buf, tag_wiretype.wire_type)\n'
				unpack_text += 'res.$name << v\n'
				unpack_text += 'i = ii\n'
				unpack_text += '}\n'
			} else {
				pack_text += '// [packed=true]\n'
				pack_text += 'res << ${pack_inside}_packed(o.$name, $number)\n'
				
				unpack_text += '$number {\n'
				unpack_text += '// [packed=true]\n'
				unpack_text += 'ii, v := ${unpack_inside}_packed(cur_buf, tag_wiretype.wire_type)\n'
				unpack_text += 'res.$name << v\n'
				unpack_text += 'i = ii\n'
				unpack_text += '}\n'
			}
		}

		else {
			// This should never happen...
			println('Unknown label $label')
		}
	}

	return pack_text, unpack_text
}

fn key_default_value(v_type string) string {
	match v_type {
		'string' {
			return '\'\''
		}

		'[]byte' {
			// Keys cant be this type but value_default_value uses this for
			// its .other case
			return '[]byte{}'
		}

		else {
			return '${v_type}(0)'
		}
	}
}

fn value_default_value(v_type string, type_type TypeType) string {
	match type_type {
		.other {
			return key_default_value(v_type)
		}

		else {
			return 'new_${v_type}()'
		}
	}
}

fn (g &Gen) gen_map_field_pack_text(
	key_proto_type, key_v_type, value_proto_type, value_v_type string,
	value_type_type TypeType, 
	name, number string
) (string, string){
	// TODO this isnt ideal

	value_v_type_no_mod := value_v_type.all_after_last('.')
	value_v_type_mod := if value_v_type.contains('.') { value_v_type.all_before_last('.') + '.' } else { '' }

	value_pack_inside := g.type_pack_name('${value_v_type_mod}pack', value_proto_type, value_v_type_no_mod, value_type_type)
	value_unpack_inside := g.type_pack_name('${value_v_type_mod}unpack', value_proto_type, value_v_type_no_mod, value_type_type)

	key_pack_inside := g.type_pack_name('pack', key_proto_type, key_v_type, .other)
	key_unpack_inside := g.type_pack_name('unpack', key_proto_type, key_v_type, .other)


	mut pack_text := ''
	mut unpack_text := ''
	// Essentially the same as a repeated field of a message
	// where the message first contains the key
	// and then the value
	pack_text += 'for k, v in o.$name {\n'
	pack_text += 'mut bytes := ${key_pack_inside}(k, 1)'
	pack_text += 'bytes << ${value_pack_inside}(v, 2)'
	pack_text += 'res << vproto.pack_bytes_field(bytes, $number)'
	pack_text += '}\n'

	unpack_text += '$number {\n'
	unpack_text += 'ii, bytes := vproto.unpack_message_field(cur_buf, tag_wiretype.wire_type)\n'
	unpack_text += 'mut k := ${key_default_value(key_v_type)}\n'
	unpack_text += 'mut v := ${value_default_value(value_v_type, value_type_type)}\n'
	unpack_text += 'mut bytes_offset := 0\n'
	unpack_text += 'for j := 0; j < 2; j++ {\n'
	unpack_text += 'map_tag_wiretype := vproto.unpack_tag_wire_type(bytes[bytes_offset..]) or { return error(\'malformed protobuf (couldnt parse tag & wire type)\') }\n'
	unpack_text += 'match map_tag_wiretype.tag {\n'
	unpack_text += '1 {\n'
	unpack_text += 'map_ii, kk := ${key_unpack_inside}(bytes[bytes_offset..],  map_tag_wiretype.wire_type)\n'
	unpack_text += 'bytes_offset += map_ii\n'
	unpack_text += 'k = kk\n'
	unpack_text += '}\n'
	unpack_text += '2 {\n'
	unpack_text += 'map_ii, vv := ${value_unpack_inside}(bytes[bytes_offset..], map_tag_wiretype.wire_type) \n'
	unpack_text += 'bytes_offset += map_ii\n'
	unpack_text += 'v = vv\n'
	unpack_text += '}\n'
	unpack_text += 'else { \n'
	unpack_text += 'return error(\'malformed map field (didnt unpack a key/value)\')\n'
	unpack_text += '}\n'
	unpack_text += '}\n'
	unpack_text += '}\n'
	unpack_text += 'res.$name[k] = v\n'
	unpack_text += 'i = ii\n'
	unpack_text += '}\n'

	return pack_text, unpack_text
}

fn (mut g Gen) gen_message_internal(type_context []string, m &Message) {
	m_names := g.message_names(type_context, m.name)

	m_name := m_names.struct_name
	m_full_name := m_names.lowercase_name

	// Generate for submessages
	for _, sub in m.messages {
		g.gen_message_internal(m_names.this_type_context, sub)
	}
	
	// Generate for subenums
	for _, sub in m.enums {
		g.gen_enum_definition(m_names.this_type_context, sub)
	}

	has_fields := 0 < m.fields.len + m.map_fields.len

	pack_unpack_mut := if has_fields {
		'mut '
	} else {
		''
	}

	mut field_pack_text := new_writer()
	mut field_unpack_text := new_writer()

	field_pack_text.l('pub fn (o &$m_name) pack() []byte {')
	field_pack_text.l('${pack_unpack_mut}res := []byte{}') // TODO allocate correct size statically
	
	field_unpack_text.l('pub fn ${m_full_name}_unpack(buf []byte) ?$m_name {')
	field_unpack_text.l('${pack_unpack_mut}res := $m_name{}')

	if has_fields {
		field_unpack_text.l('mut total := 0')
		field_unpack_text.l('for total < buf.len {')
		field_unpack_text.l('mut i := 0')
		field_unpack_text.l('buf_before_wire_type := buf[total..]')
		field_unpack_text.l('tag_wiretype := vproto.unpack_tag_wire_type(buf_before_wire_type) or { return error(\'malformed protobuf (couldnt parse tag & wire type)\') }')
		field_unpack_text.l('cur_buf := buf_before_wire_type[tag_wiretype.consumed..]')
		field_unpack_text.l('match tag_wiretype.tag {')
	}

	g.w.l('pub struct $m_name {')

	g.w.l('mut:')
	g.w.l('unknown_fields []vproto.UnknownField')


	if has_fields {
		g.w.l('pub mut:')
	}

	for field in m.fields {
		// simple_context := simplify_type_context(field.type_context, type_context)
		// println('$type_context - $field.type_context = $simple_context')
		field_type, field_type_type := g.type_to_typename(field.type_context, field.t)

		name := escape_name(field.name)

		if field.label == 'optional' {
			g.w.l('${name} ${field_type}')
			g.w.l('has_${name} bool')

		} else if field.label == 'required' {
			g.w.l('${name} ${field_type}')
		} else if field.label == 'repeated' {
			g.w.l('${name} []${field_type}')
		}

		mut is_packed := false
		if field.label == 'repeated' {
			for o in field.options {
				if o.ident == 'packed' {
					is_packed = o.value.value == 'true'
				}
			}
		}

		mut pack_text := ''
		mut unpack_text := ''

		if field_type_type == .enum_ || field_type_type == .message {
			names := g.message_names(field.type_context, field.t)

			// n := (field.type_context.join('') + names.lowercase_name).to_lower()
			pack_text, unpack_text = g.gen_field_pack_text(field.label, field.t, names.lowercase_name, field_type_type, name, field.number, is_packed)
		} else {
			pack_text, unpack_text = g.gen_field_pack_text(field.label, field.t, field_type, field_type_type, name, field.number, is_packed)
		}

		field_pack_text.l(pack_text)
		field_unpack_text.l(unpack_text)
	}

	for map_field in m.map_fields {
		key_type, _ := g.type_to_typename(map_field.type_context, map_field.key_type)
		value_type, value_type_type := g.type_to_typename(map_field.type_context, map_field.value_type)

		name := escape_name(map_field.name)

		g.w.l('${name} map[$key_type]$value_type')

		mut pack_text := ''
		mut unpack_text := ''

		if value_type_type == .enum_ || value_type_type == .message {
			names := g.message_names(map_field.type_context, map_field.value_type)

			pack_text, unpack_text = g.gen_map_field_pack_text(map_field.key_type, key_type, map_field.value_type, names.lowercase_name, value_type_type, name, map_field.number)
		} else {
			pack_text, unpack_text = g.gen_map_field_pack_text(map_field.key_type, key_type, map_field.value_type, value_type, value_type_type, name, map_field.number)
		}

		field_pack_text.l(pack_text)
		field_unpack_text.l(unpack_text)
	}

	// TODO oneofs maps extensions and similar

	g.w.l('}')

	field_pack_text.l('return res')
	field_pack_text.l('}')

	if has_fields {
		// close match then for then func
		field_unpack_text.l('else {')
		field_unpack_text.l('ii, v := vproto.unpack_unknown_field(cur_buf, tag_wiretype.wire_type)')
		field_unpack_text.l('res.unknown_fields << vproto.UnknownField{tag_wiretype.wire_type, tag_wiretype.tag, v}')
		field_unpack_text.l('i = ii')
		field_unpack_text.l('}')
		field_unpack_text.l('}')

		// TODO we need to actually implement parsing of unknown fields otherwise this will
		// always trigger if we hit one
		field_unpack_text.l('if i == 0 { return error(\'malformed protobuf (didnt unpack a field)\') }')
		field_unpack_text.l('total += tag_wiretype.consumed + i')
		field_unpack_text.l('}')
	}
	field_unpack_text.l('return res')
	field_unpack_text.l('}')

	// Function for creating a new of that message

	g.w.l('pub fn new_${m_full_name}() $m_name {')
	g.w.l('return $m_name{}')
	g.w.l('}')

	g.w.l(field_pack_text.text())
	g.w.l(field_unpack_text.text())

	// pack and unpack wrappers for when its called as a submessage
	g.w.l('pub fn pack_${m_full_name}(o $m_name, num u32) []byte {')
	g.w.l('return vproto.pack_message_field(o.pack(), num)')
	g.w.l('}')
	
	g.w.l('pub fn unpack_${m_full_name}(buf []byte, tag_wiretype vproto.WireType) (int, $m_name) {')
	g.w.l('i, v := vproto.unpack_message_field(buf, tag_wiretype)')
	g.w.l('unpacked := ${m_full_name}_unpack(v) or { panic(\'\') }')
	g.w.l('return i, unpacked')
	g.w.l('}')

	// TODO oneof, maps and similar
}

pub fn (mut g Gen) gen_file_text(f &File) string {
	g.current_package = f.package
	g.gen_file_header(f)

	for _, e in f.enums {
		g.gen_enum_definition([f.package], e)
	}

	// Then generate the actual structs that back the messages
	for _, m in f.messages {
		g.gen_message_internal([f.package], m)
	}

	return g.w.text()
}

pub fn new_gen(p &Parser) Gen {
	mut g := Gen{type_table: p.type_table, w: new_writer()}

	for _, f in p.files {
		mod := f.package

		g.package_lookup[f.filename] = mod
	}

	return g
}